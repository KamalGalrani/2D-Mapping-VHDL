library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity D_Lookup is
  port(
      THETA2 : in  integer range -360 to 360;
      DX     : out integer range -15 to 15;
      DY     : out integer range -15 to 15;
      DT     : out integer range 0 to 7
      );
end entity;

architecture main of D_Lookup is
signal theta2_a         : integer range 0 to 360;
signal theta2_r         : integer range 0 to 180;
signal neg_dx, neg_dy   : std_logic := '0';
signal dx_buff, dy_buff : integer range 0 to 15;
begin
  DT <= 1;
  theta2_r <= abs(THETA2) when ( abs(THETA2) <= 180 )
                      else 360 - abs(THETA2);

  DY       <= dy_buff     when ( abs(THETA2) <= 180 )
                      else -1*dy_buff;

  DX       <= dx_buff      when ( THETA2 >= 0 )
                      else -1*dx_buff;

with theta2_r select
dy_buff <=  0 when 180,
            0 when 179,
            0 when 178,
            0 when 177,
            0 when 176,
            0 when 175,
            0 when 174,
            1 when 173,
            1 when 172,
            1 when 171,
            1 when 170,
            1 when 169,
            1 when 168,
            1 when 167,
            1 when 166,
            1 when 165,
            1 when 164,
            1 when 163,
            1 when 162,
            1 when 161,
            2 when 160,
            2 when 159,
            2 when 158,
            2 when 157,
            2 when 156,
            2 when 155,
            2 when 154,
            2 when 153,
            2 when 152,
            2 when 151,
            2 when 150,
            2 when 149,
            2 when 148,
            2 when 147,
            3 when 146,
            3 when 145,
            3 when 144,
            3 when 143,
            3 when 142,
            3 when 141,
            3 when 140,
            3 when 139,
            3 when 138,
            3 when 137,
            3 when 136,
            3 when 135,
            3 when 134,
            3 when 133,
            4 when 132,
            4 when 131,
            4 when 130,
            4 when 129,
            4 when 128,
            4 when 127,
            4 when 126,
            4 when 125,
            4 when 124,
            4 when 123,
            4 when 122,
            4 when 121,
            4 when 120,
            4 when 119,
            4 when 118,
            5 when 117,
            5 when 116,
            5 when 115,
            5 when 114,
            5 when 113,
            5 when 112,
            5 when 111,
            5 when 110,
            5 when 109,
            5 when 108,
            5 when 107,
            5 when 106,
            5 when 105,
            5 when 104,
            5 when 103,
            5 when 102,
            6 when 101,
            6 when 100,
            6 when 99,
            6 when 98,
            6 when 97,
            6 when 96,
            6 when 95,
            6 when 94,
            6 when 93,
            6 when 92,
            6 when 91,
            6 when 90,
            6 when 89,
            6 when 88,
            6 when 87,
            6 when 86,
            6 when 85,
            6 when 84,
            7 when 83,
            7 when 82,
            7 when 81,
            7 when 80,
            7 when 79,
            7 when 78,
            7 when 77,
            7 when 76,
            7 when 75,
            7 when 74,
            7 when 73,
            7 when 72,
            7 when 71,
            7 when 70,
            7 when 69,
            7 when 68,
            7 when 67,
            7 when 66,
            7 when 65,
            7 when 64,
            7 when 63,
            7 when 62,
            8 when 61,
            8 when 60,
            8 when 59,
            8 when 58,
            8 when 57,
            8 when 56,
            8 when 55,
            8 when 54,
            8 when 53,
            8 when 52,
            8 when 51,
            8 when 50,
            8 when 49,
            8 when 48,
            8 when 47,
            8 when 46,
            8 when 45,
            8 when 44,
            8 when 43,
            8 when 42,
            8 when 41,
            8 when 40,
            8 when 39,
            8 when 38,
            8 when 37,
            8 when 36,
            8 when 35,
            8 when 34,
            8 when 33,
            8 when 32,
            8 when 31,
            8 when 30,
            8 when 29,
            8 when 28,
            8 when 27,
            9 when 26,
            9 when 25,
            9 when 24,
            9 when 23,
            9 when 22,
            9 when 21,
            9 when 20,
            9 when 19,
            9 when 18,
            9 when 17,
            9 when 16,
            9 when 15,
            9 when 14,
            9 when 13,
            9 when 12,
            9 when 11,
            9 when 10,
            9 when 9,
            9 when 8,
            9 when 7,
            9 when 6,
            9 when 5,
            9 when 4,
            9 when 3,
            9 when 2,
            9 when 1,
            9 when 0,
            9 when others;

with theta2_r select
dx_buff <=  0 when 0,
            0 when 1,
            0 when 2,
            0 when 3,
            0 when 4,
            0 when 5,
            0 when 6,
            1 when 7,
            1 when 8,
            1 when 9,
            1 when 10,
            1 when 11,
            1 when 12,
            1 when 13,
            1 when 14,
            1 when 15,
            1 when 16,
            1 when 17,
            1 when 18,
            1 when 19,
            2 when 20,
            2 when 21,
            2 when 22,
            2 when 23,
            2 when 24,
            2 when 25,
            2 when 26,
            2 when 27,
            2 when 28,
            2 when 29,
            2 when 30,
            2 when 31,
            2 when 32,
            2 when 33,
            3 when 34,
            3 when 35,
            3 when 36,
            3 when 37,
            3 when 38,
            3 when 39,
            3 when 40,
            3 when 41,
            3 when 42,
            3 when 43,
            3 when 44,
            3 when 45,
            3 when 46,
            3 when 47,
            4 when 48,
            4 when 49,
            4 when 50,
            4 when 51,
            4 when 52,
            4 when 53,
            4 when 54,
            4 when 55,
            4 when 56,
            4 when 57,
            4 when 58,
            4 when 59,
            4 when 60,
            4 when 61,
            4 when 62,
            5 when 63,
            5 when 64,
            5 when 65,
            5 when 66,
            5 when 67,
            5 when 68,
            5 when 69,
            5 when 70,
            5 when 71,
            5 when 72,
            5 when 73,
            5 when 74,
            5 when 75,
            5 when 76,
            5 when 77,
            5 when 78,
            6 when 79,
            6 when 80,
            6 when 81,
            6 when 82,
            6 when 83,
            6 when 84,
            6 when 85,
            6 when 86,
            6 when 87,
            6 when 88,
            6 when 89,
            6 when 90,
            6 when 91,
            6 when 92,
            6 when 93,
            6 when 94,
            6 when 95,
            6 when 96,
            7 when 97,
            7 when 98,
            7 when 99,
            7 when 100,
            7 when 101,
            7 when 102,
            7 when 103,
            7 when 104,
            7 when 105,
            7 when 106,
            7 when 107,
            7 when 108,
            7 when 109,
            7 when 110,
            7 when 111,
            7 when 112,
            7 when 113,
            7 when 114,
            7 when 115,
            7 when 116,
            7 when 117,
            7 when 118,
            8 when 119,
            8 when 120,
            8 when 121,
            8 when 122,
            8 when 123,
            8 when 124,
            8 when 125,
            8 when 126,
            8 when 127,
            8 when 128,
            8 when 129,
            8 when 130,
            8 when 131,
            8 when 132,
            8 when 133,
            8 when 134,
            8 when 135,
            8 when 136,
            8 when 137,
            8 when 138,
            8 when 139,
            8 when 140,
            8 when 141,
            8 when 142,
            8 when 143,
            8 when 144,
            8 when 145,
            8 when 146,
            8 when 147,
            8 when 148,
            8 when 149,
            8 when 150,
            8 when 151,
            8 when 152,
            8 when 153,
            9 when 154,
            9 when 155,
            9 when 156,
            9 when 157,
            9 when 158,
            9 when 159,
            9 when 160,
            9 when 161,
            9 when 162,
            9 when 163,
            9 when 164,
            9 when 165,
            9 when 166,
            9 when 167,
            9 when 168,
            9 when 169,
            9 when 170,
            9 when 171,
            9 when 172,
            9 when 173,
            9 when 174,
            9 when 175,
            9 when 176,
            9 when 177,
            9 when 178,
            9 when 179,
            9 when 180,
            0 when others;

end architecture;
