library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity UART is
  generic(
		-------------------------------------------------
      --TX_CLK_DIV = FCPU/BAUDRATE - 1
        --9600   => 5207
        --14400  => 3471
        --19200  => 2603
        --28800  => 1735
        --38400  => 1301
        --57600  => 867
        --115200 => 433
      -------------------------------------------------
      TX_CLK_DIV : integer := 5207
      );
  port(
      CLK   : in  std_logic;
      RST   : in  std_logic;
      WR    : in  std_logic;
      TX    : out std_logic;
      TXRDY : out std_logic
      );
end entity;

architecture main of UART is
signal tx_clk_count : integer range 0 to TX_CLK_DIV;
signal tx_clk_tick  : std_logic;
signal TX_DATA: std_logic_vector(7 downto 0);
component TRANSMIT is
  port(
      TX_CLK : in std_logic;
      WR     : in std_logic;
      RST    : in std_logic;
      DATA   : in std_logic_vector(7 downto 0);
      TX     : out std_logic;
      TXRDY  : out std_logic
		);
end component;
begin
  process (RST, CLK)
  begin
    if ( RST = '1' ) then
      tx_clk_tick  <= '0';
      tx_clk_count <= 0;
    elsif rising_edge(CLK) then
      tx_clk_tick <= '0';
      if (tx_clk_count = TX_CLK_DIV) then
        tx_clk_count <= 0;
        tx_clk_tick <= '1';
      else
        tx_clk_count <= tx_clk_count + 1;
      end if;
    end if;
  end process;
  transmitter: TRANSMIT port map (tx_clk_tick, WR, RST, "01000010", TX, TXRDY);
end architecture;