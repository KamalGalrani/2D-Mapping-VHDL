library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ADC is 
  port(
      ADC  : in  unsigned(7 downto 0);
		DIST : out integer range 0 to 1300
      );
end entity;

architecture main of ADC is
begin
  with to_integer(ADC) select
    DIST <= 0 when 255,
            5 when 254,
            10 when 253,
            15 when 252,
            20 when 251,
            25 when 250,
            30 when 249,
            35 when 248,
            40 when 247,
            45 when 246,
            50 when 245,
            56 when 244,
            61 when 243,
            66 when 242,
            71 when 241,
            76 when 240,
            81 when 239,
            86 when 238,
            91 when 237,
            96 when 236,
            101 when 235,
            107 when 234,
            112 when 233,
            117 when 232,
            122 when 231,
            127 when 230,
            132 when 229,
            137 when 228,
            142 when 227,
            147 when 226,
            152 when 225,
            158 when 224,
            163 when 223,
            168 when 222,
            173 when 221,
            178 when 220,
            183 when 219,
            188 when 218,
            193 when 217,
            198 when 216,
            203 when 215,
            209 when 214,
            214 when 213,
            219 when 212,
            224 when 211,
            229 when 210,
            234 when 209,
            239 when 208,
            244 when 207,
            249 when 206,
            254 when 205,
            260 when 204,
            265 when 203,
            270 when 202,
            275 when 201,
            280 when 200,
            285 when 199,
            290 when 198,
            295 when 197,
            300 when 196,
            305 when 195,
            310 when 194,
            316 when 193,
            321 when 192,
            326 when 191,
            331 when 190,
            336 when 189,
            341 when 188,
            346 when 187,
            351 when 186,
            356 when 185,
            361 when 184,
            367 when 183,
            372 when 182,
            377 when 181,
            382 when 180,
            387 when 179,
            392 when 178,
            397 when 177,
            402 when 176,
            407 when 175,
            412 when 174,
            418 when 173,
            423 when 172,
            428 when 171,
            433 when 170,
            438 when 169,
            443 when 168,
            448 when 167,
            453 when 166,
            458 when 165,
            463 when 164,
            469 when 163,
            474 when 162,
            479 when 161,
            484 when 160,
            489 when 159,
            494 when 158,
            499 when 157,
            504 when 156,
            509 when 155,
            514 when 154,
            520 when 153,
            525 when 152,
            530 when 151,
            535 when 150,
            540 when 149,
            545 when 148,
            550 when 147,
            555 when 146,
            560 when 145,
            565 when 144,
            570 when 143,
            576 when 142,
            581 when 141,
            586 when 140,
            591 when 139,
            596 when 138,
            601 when 137,
            606 when 136,
            611 when 135,
            616 when 134,
            621 when 133,
            627 when 132,
            632 when 131,
            637 when 130,
            642 when 129,
            647 when 128,
            652 when 127,
            657 when 126,
            662 when 125,
            667 when 124,
            672 when 123,
            678 when 122,
            683 when 121,
            688 when 120,
            693 when 119,
            698 when 118,
            703 when 117,
            708 when 116,
            713 when 115,
            718 when 114,
            723 when 113,
            729 when 112,
            734 when 111,
            739 when 110,
            744 when 109,
            749 when 108,
            754 when 107,
            759 when 106,
            764 when 105,
            769 when 104,
            774 when 103,
            780 when 102,
            785 when 101,
            790 when 100,
            795 when 99,
            800 when 98,
            805 when 97,
            810 when 96,
            815 when 95,
            820 when 94,
            825 when 93,
            830 when 92,
            836 when 91,
            841 when 90,
            846 when 89,
            851 when 88,
            856 when 87,
            861 when 86,
            866 when 85,
            871 when 84,
            876 when 83,
            881 when 82,
            887 when 81,
            892 when 80,
            897 when 79,
            902 when 78,
            907 when 77,
            912 when 76,
            917 when 75,
            922 when 74,
            927 when 73,
            932 when 72,
            938 when 71,
            943 when 70,
            948 when 69,
            953 when 68,
            958 when 67,
            963 when 66,
            968 when 65,
            973 when 64,
            978 when 63,
            983 when 62,
            989 when 61,
            994 when 60,
            999 when 59,
            1004 when 58,
            1009 when 57,
            1014 when 56,
            1019 when 55,
            1024 when 54,
            1029 when 53,
            1034 when 52,
            1040 when 51,
            1045 when 50,
            1050 when 49,
            1055 when 48,
            1060 when 47,
            1065 when 46,
            1070 when 45,
            1075 when 44,
            1080 when 43,
            1085 when 42,
            1090 when 41,
            1096 when 40,
            1101 when 39,
            1106 when 38,
            1111 when 37,
            1116 when 36,
            1121 when 35,
            1126 when 34,
            1131 when 33,
            1136 when 32,
            1141 when 31,
            1147 when 30,
            1152 when 29,
            1157 when 28,
            1162 when 27,
            1167 when 26,
            1172 when 25,
            1177 when 24,
            1182 when 23,
            1187 when 22,
            1192 when 21,
            1198 when 20,
            1203 when 19,
            1208 when 18,
            1213 when 17,
            1218 when 16,
            1223 when 15,
            1228 when 14,
            1233 when 13,
            1238 when 12,
            1243 when 11,
            1249 when 10,
            1254 when 9,
            1259 when 8,
            1264 when 7,
            1269 when 6,
            1274 when 5,
            1279 when 4,
            1284 when 3,
            1289 when 2,
            1294 when 1,
            1300 when 0,
				0    when others;
end architecture;